-- Code your design here
-- Code your design here
library IEEE;
use IEEE.std_logic_1164.all;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

Entity Buffers is
port (
	clk : in std_logic;
    reset : in std_logic;
	Mem1_in : in std_logic_vector(7 downto 0);
    Mem1_out : out std_logic_vector(7 downto 0);
    MEM1_val : in std_logic;
    
    Mem2_in : in std_logic_vector(7 downto 0);
    Mem2_out : in std_logic_vector(7 downto 0);
    Mem2_val : in std_logic;
    
    SR_L_in : in std_logic;
    SR_L_in : in std_logic;
    SR_L_val : in std_logic;
    
    SR_R_out : in std_logic;
    SR_R_out : in std_logic;
    SR_L_val : in std_logic;
    
    BuffA_in : in std_logic_vector(3 downto 0);
    BuffA_out : in std_logic_vector(3 downto 0);
    BuffA_val : std_logic;
    
    BuffB_in : in std_logic_vector(3 downto 0);
    BuffB_out : in std_logic_vector(3 downto 0);
    BuffB_val : std_logic;
  	)
    end Buffers;
architecture Buffers_arch of Buffers is
begin
	BuffA_process : process (reset,clk,BuffA_val)
    begin 
 		if reset ='1' then
        	BuffA_out <= (other => '0');
        else if (rising_edge (clk) and BuffA_val ='0') then
        	BuffA_out <= BuffA_in;
    	end if;
    end process;